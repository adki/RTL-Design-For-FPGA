//--------------------------------------------------------
// Copyright (c) 2020 by Ando Ki.
// All right reserved.
//
// http://www.future-ds.com
// adki@future-ds.com
//--------------------------------------------------------
`timescale 1ns/1ns

module top ;
   //--------------------------------------------------------
   ...
   //--------------------------------------------------------
   apb_gpio_tester u_tester (
      .........
   );
   //--------------------------------------------------------
   gpio_apb #(.GPIO_WIDTH(GPIO_WIDTH))
   u_gpio (
       ............
   );
endmodule
