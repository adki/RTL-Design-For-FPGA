/**********************************************************
Proxy module for full_adder
Generated automatically by iNSPIRE at  12:58:34 02/21/09
**********************************************************/
module full_adder (
  clk,
  cout,
  sum,
  resetb,
  in1,
  in2,
  cin  );

  input clk;
  output cout;
  output sum;
  input resetb;
  input in1;
  input in2;
  input cin;

  reg cout;
  reg sum;
  // Internal nodes


  initial $iProveEmulation;

endmodule
