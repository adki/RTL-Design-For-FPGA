/*
 * Copyright (c) 2020 by Ando Ki.
 * All right reserved.
 *
 * http://www.future-ds.com
 * adki@future-ds.com
 *
 */
`timescale 1ns/1ns

module apb_gpio_tester (
       ...
);
   `include "apb_tasks.v"
    .............
endmodule
